// RS-�������
module RStrigger (out,x,xdop);
   // ����������� ������� � �������� ����������:
   // - x - S;
   // - xdop - R;
   // - out - !Q.
   input x,xdop;
   output out;

   // ����������� ����������� ����������
   reg res;

   // module RStrigger � �������� � RS-�������� �� �-��, � RS-�������� �� ���-��.
   // ��������������, ��� �� ������ ������ �� ��� RS-�������� ��������� ���������� ��������.
   // ��������� �������� ��������, ���� ��������� �������� ���������� x ��� xdop.
   always @(xdop or x)
   begin
      // ���� �������� �� ��������������� ������ �� ����� R, �� � ������� ����� 0
      if (~xdop)
         res = 0;
      // � ���� �������� �� ��������������� ������ �� ����� S, �� � ������� ����� 1
      else if (~x)
         res = 1;
      end
   // ����������� � ������ �������� �������� �� �����:
   assign out = !res;
endmodule

// ���������� ������
module Filter (OutResult, X, A, B);
   // ����������� ������� � �������� ����������:
   // - X - ����������� ������;
   // - A, B - �������������� �������.
   input   X, A, B;

   // �������� ���� - ��������� - ��������������� ������
   output  OutResult;

   // �������� ����������� ������, ����������� ���������� ��������
   // �������������� � ������� NOT1 � NOT2
   // ����������� ���������� � � � � ����������� ��������
   // ���������� AInv � BInv ��������������
   not NOT1 (AInv, A);
   not NOT2 (BInv, B);

   // �������� 4 ���� ������ RSTrigger, �.�. � ��� � ����� 4 ��������,
   // ���������� ��������������� ��������� ������� �������� ������� ������
   RStrigger call1 (ou1, X, A);
   RStrigger call2 (ou2, X, B);
   RStrigger call3 (ou3, X, AInv);
   RStrigger call4 (ou4, X, BInv);

   // ����� ������, ������������ ���������� �������� � � ������ AND1:
   and  AND1 (OutResult,ou1, ou2, ou3, ou4);
endmodule

