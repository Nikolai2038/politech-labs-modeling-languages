--*************************************************************
--* This file is automatically generated test bench template  *
--* By ACTIVE-VHDL    <TBgen v1.10>. Copyright (C) ALDEC Inc. *
--*                                                           *
--* This file was generated on:             20:53, 01.03.2024 *
--* Tested entity name:                                ALU_32 *
--* File name contains tested entity:        .\src\alu_32.vhd *
--*************************************************************

library ieee;
use work.dp32_types.all;
use work.alu_32_types.all;
use ieee.std_logic_1164.all;

-- Add your library and packages declaration here ...

entity alu_32_tb is
    -- Generic declarations of the tested unit
    generic (
        TPD : time := 1.0 ns
    );
end alu_32_tb;

architecture TB_ARCHITECTURE of alu_32_tb is
    -- Component declaration of the tested unit
    component ALU_32
        generic (
            TPD : time := 1.0 ns
        );
        port (
            operand1 : in bit_32;
            operand2 : in bit_32;
            result : out bus_bit_32;
            cond_code : out CC_bits;
            command : in ALU_command
        );
    end component;

    -- Stimulus signals - signals mapped to the input and inout ports of tested entity
    signal operand1 : bit_32;
    signal operand2 : bit_32;
    signal command : ALU_command;
    -- Observed signals - signals mapped to the output ports of tested entity
    signal result : bus_bit_32;
    signal cond_code : CC_bits;

    -- Add your code here ...

begin

    -- Unit Under Test port map
    UUT : ALU_32
    port map(
        operand1 => operand1,
        operand2 => operand2,
        result => result,
        cond_code => cond_code,
        command => command);

    --Below VHDL code is an inserted .\Generic\by_hand.vhs
    --User can modify it ....

    STIMULUS : process
    begin -- of stimulus process
        --wait for <time to next event>; -- <current time>

        operand2 <= "00000000000000000000000000000101";
        operand1 <= "00000000000000000000000000001011";
        command <= disable;
        wait for 100 ns; --0 ps
        command <= pass1;
        wait for 100 ns; --100 ns
        command <= log_and;
        wait for 100 ns; --200 ns
        command <= log_or;
        wait for 100 ns; --300 ns
        command <= log_xor;
        wait for 100 ns; --400 ns
        command <= log_mask;
        wait for 100 ns; --500 ns
        command <= incr1;
        wait for 100 ns; --600 ns
        command <= add;
        wait for 100 ns; --700 ns
        command <= subtract;
        wait for 100 ns; --800 ns
        command <= multiply;
        wait for 100 ns; --900 ns
        --    end of stimulus events
        wait;
    end process; -- end of stimulus process

    -- Add your stimulus here ...

end TB_ARCHITECTURE;

configuration TESTBENCH_FOR_ALU_32 of alu_32_tb is
    for TB_ARCHITECTURE
        for UUT : ALU_32
            use entity work.ALU_32(behaviour);
        end for;
    end for;
end TESTBENCH_FOR_ALU_32;
