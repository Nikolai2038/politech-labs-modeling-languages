--*************************************************************
--* This file is automatically generated test bench template  *
--* By ACTIVE-VHDL    <TBgen v1.10>. Copyright (C) ALDEC Inc. *
--*                                                           *
--* This file was generated on:              2:33, 20.05.2024 *
--* Tested entity name:                                  sort *
--* File name contains tested entity:          .\src\sort.vhd *
--*************************************************************

library ieee;
use work.sort_types.all;
use ieee.std_logic_1164.all;

	-- Add your library and packages declaration here ...

entity sort_tb is
end sort_tb;

architecture TB_ARCHITECTURE of sort_tb is
	-- Component declaration of the tested unit
	component sort
	port(
		clk : in std_logic;
		reset : in std_logic;
		working : out std_logic;
		data_in : in massType;
		data_out : out massType );
end component;

	-- Stimulus signals - signals mapped to the input and inout ports of tested entity
	signal clk : std_logic;
	signal reset : std_logic;
	signal data_in : massType;
	-- Observed signals - signals mapped to the output ports of tested entity
	signal working : std_logic;
	signal data_out : massType;

	-- Add your code here ...

begin

	-- Unit Under Test port map
	UUT : sort
		port map
			(clk => clk,
			reset => reset,
			working => working,
			data_in => data_in,
			data_out => data_out );

	--Below VHDL code is an inserted .\Generic\sort_waveform.vhs
	--User can modify it ....

STIMULUS: process
begin  -- of stimulus process
--wait for <time to next event>; -- <current time>

--	end of stimulus events
	wait;
end process; -- end of stimulus process
	



	-- Add your stimulus here ...

end TB_ARCHITECTURE;

configuration TESTBENCH_FOR_sort of sort_tb is
	for TB_ARCHITECTURE
		for UUT : sort
			use entity work.sort(sort_architecture);
		end for;
	end for;
end TESTBENCH_FOR_sort;

